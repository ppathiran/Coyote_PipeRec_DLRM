always_comb begin 
    /*
     * CONTROL SIGNALS
     * 
     * rq_(wr|rd) are two more Coyote interfaces, which act as inputs to the user application
     * They corresponds to network write/read requests, set from the host software and driver
     * Here, they are used to set Coyote's generic send queues, previously discussed in Example 7.
     */
    // Write
    sq_wr.valid = rq_wr.valid;
    rq_wr.ready = sq_wr.ready;
    sq_wr.data = rq_wr.data;            // Data field holds information such as remote, virtual address, buffer length etc.
    sq_wr.data.strm = STRM_HOST;        // For RDMA, by definition data is always on the host
    sq_wr.data.dest = is_opcode_rd_resp(rq_wr.data.opcode) ? 0 : 1;

    // Reads
    sq_rd.valid = rq_rd.valid;
    rq_rd.ready = sq_rd.ready;
    sq_rd.data = rq_rd.data;           // Data field holds information such as remote, virtual address, buffer length etc.
    sq_rd.data.strm = STRM_HOST;       // For RDMA, by definition data is always on the host
    sq_rd.data.dest = 1;
end

/*
 * DATA SIGNALS
 * 
 */


// Data streams for outgoing RDMA WRITEs (from local host to network stack to remote node)
`AXISR_ASSIGN(axis_host_recv[0], axis_rreq_send[0])

// Data streams for incoming RDMA READ RESPONSEs (from remote node to network stack to local host)
// `AXISR_ASSIGN(axis_rreq_recv[0], axis_host_send[0])


hls_vadd inst_vadd(
    .s_axi_in_TDATA        (axis_rreq_recv[0].tdata),
    .s_axi_in_TKEEP        (axis_rreq_recv[0].tkeep),
    .s_axi_in_TLAST        (axis_rreq_recv[0].tlast),
    .s_axi_in_TSTRB        (0),
    .s_axi_in_TVALID       (axis_rreq_recv[0].tvalid),
    .s_axi_in_TREADY       (axis_rreq_recv[0].tready),

    .m_axi_out_TDATA        (axis_host_send[0].tdata),
    .m_axi_out_TKEEP        (axis_host_send[0].tkeep),
    .m_axi_out_TLAST        (axis_host_send[0].tlast),
    .m_axi_out_TSTRB        (),
    .m_axi_out_TVALID       (axis_host_send[0].tvalid),
    .m_axi_out_TREADY       (axis_host_send[0].tready),

    .ap_clk                 (aclk),
    .ap_rst_n               (aresetn)
);


// Data streams for outgoing RDMA READ RESPONSEs (from local host to network stack to remote node)
`AXISR_ASSIGN(axis_host_recv[1], axis_rrsp_send[0])

// Data streams for incoming RDMA WRITEs (from remote node to network stack to local host)
`AXISR_ASSIGN(axis_rrsp_recv[0], axis_host_send[1])

// Tie off unused interfaces
always_comb axi_ctrl.tie_off_s();
always_comb notify.tie_off_m();
always_comb cq_rd.tie_off_s();
always_comb cq_wr.tie_off_s();

// // ILA for debugging
// ila_perf_rdma inst_ila_perf_rdma (
//     .clk(aclk),
//     .probe0(axis_host_recv[0].tvalid),      // 1
//     .probe1(axis_host_recv[0].tready),      // 1
//     .probe2(axis_host_recv[0].tlast),       // 1

//     .probe3(axis_host_recv[1].tvalid),      // 1
//     .probe4(axis_host_recv[1].tready),      // 1
//     .probe5(axis_host_recv[1].tlast),       // 1

//     .probe6(axis_host_send[0].tvalid),      // 1
//     .probe7(axis_host_send[0].tready),      // 1
//     .probe8(axis_host_send[0].tlast),       // 1

//     .probe9(axis_host_send[1].tvalid),      // 1
//     .probe10(axis_host_send[1].tready),     // 1
//     .probe11(axis_host_send[1].tlast),      // 1

//     .probe12(sq_wr.valid),                  // 1
//     .probe13(sq_wr.ready),                  // 1
//     .probe14(sq_wr.data),                   // 128
//     .probe15(sq_rd.valid),                  // 1
//     .probe16(sq_rd.ready),                  // 1
//     .probe17(sq_rd.data)                    // 128
// );
